//------------------------------------------------------------------------------
// Company: 		 UIUC ECE Dept.
// Engineer:		 Stephen Kempf
//
// Create Date:    
// Design Name:    ECE 385 Lab 5 Given Code - SLC-3 top-level (Physical RAM)
// Module Name:    SLC3
//
// Comments:
//    Revised 03-22-2007
//    Spring 2007 Distribution
//    Revised 07-26-2013
//    Spring 2015 Distribution
//    Revised 09-22-2015 
//    Revised 06-09-2020
//	  Revised 03-02-2021
//------------------------------------------------------------------------------


module slc3(
	input logic [9:0] SW,
	input logic	Clk, Reset, Run, Continue,
	output logic [9:0] LED,
	input logic [15:0] Data_from_SRAM,
	output logic OE, WE,
	output logic [6:0] HEX0, HEX1, HEX2, HEX3,
	output logic [15:0] ADDR,
	output logic [15:0] Data_to_SRAM
);


// An array of 4-bit wires to connect the hex_drivers efficiently to wherever we want
// For Lab 1, they will direclty be connected to the IR register through an always_comb circuit
// For Lab 2, they will be patched into the MEM2IO module so that Memory-mapped IO can take place
logic [3:0] hex_4[3:0]; 
HexDriver hex_drivers[3:0] (hex_4, {HEX3, HEX2, HEX1, HEX0});
// This works thanks to http://stackoverflow.com/questions/1378159/verilog-can-we-have-an-array-of-custom-modules




// Internal connections
logic LD_MAR, LD_MDR, LD_IR, LD_BEN, LD_CC, LD_REG, LD_PC, LD_LED;
logic GatePC, GateMDR, GateALU, GateMARMUX;
logic SR2MUX, ADDR1MUX, MARMUX;
logic BEN, MIO_EN, DRMUX, SR1MUX;
logic [1:0] PCMUX, ADDR2MUX, ALUK;
logic [15:0] MDR_In;
logic [15:0] MAR, MDR, IR, PC;
logic [15:0] SR1OUT, SR2OUT, SR2MUXOUT, ADDR1MUXOUT, ADDR2MUXOUT, ALUOut, ADDRAdd;
logic [2:0] SR1MUXOUT, DRMUXOUT, CC;
logic [15:0] databus, newPC, newMDR;
logic [2:0] newCC;
logic newBEN;
logic [15:0] IR40SEXT, IR50SEXT, IR80SEXT, IR100SEXT;

//assign LED[0] = Run; 
//assign LED[1] = Continue; 
assign LED[9:0] = IR[9:0];

// Connect MAR to ADDR, which is also connected as an input into MEM2IO
//	MEM2IO will determine what gets put onto Data_CPU (which serves as a potential
//	input into MDR)
assign ADDR = MAR; 
assign MIO_EN = OE;
assign newCC = databus[15] ? 3'b100 : ((databus == 16'h0000) ? 3'b010 : 3'b001);
assign newBEN = (IR[11] & CC[2]) || (IR[10] & CC[1]) || (IR[9] & CC[0]);
assign IR40SEXT = IR[4] ? {11'hFFF, IR[4:0]} : {11'h000, IR[4:0]};
assign IR50SEXT = IR[5] ? {10'hFFF, IR[5:0]} : {10'h000, IR[5:0]};
assign IR80SEXT = IR[8] ? {7'hFF, IR[8:0]} : {7'h00, IR[8:0]};
assign IR100SEXT = IR[10] ? {5'b11111, IR[10:0]} : {5'b00000, IR[10:0]};
assign ADDRAdd = ADDR1MUXOUT + ADDR2MUXOUT;
// Connect everything to the data path (you have to figure out this part)
datapath d0 (.*);

mux_2_1 MDRMux(.in0(databus), .in1(MDR_In), .select(MIO_EN), .out(newMDR));
mux_3_1 PCMux(.in0(PC + 16'h0001), .in1(databus), .in2(ADDRAdd), .select(PCMUX), .out(newPC));
mux_2_1 #(3) SR1mux(.in0(IR[11:9]), .in1(IR[8:6]), .select(SR1MUX), .out(SR1MUXOUT));
mux_2_1 #(3) DRmux(.in0(IR[11:9]), .in1(3'b111), .select(DRMUX), .out(DRMUXOUT));
mux_2_1 SR2mux(.in0(SR2OUT), .in1(IR40SEXT), .select(SR2MUX), .out(SR2MUXOUT));
mux_2_1 ADDR1mux(.in0(PC), .in1(SR1OUT), .select(ADDR1MUX), .out(ADDR1MUXOUT));
mux_4_1 ADDR2mux(.in0(16'h0000), .in1(IR50SEXT), .in2(IR80SEXT), .in3(IR100SEXT), .select(ADDR2MUX), .out(ADDR2MUXOUT));
fetch_reg_unit fetch(.*, .PCIn(newPC), .MARIn(databus), .MDRIn(newMDR), .IRIn(databus), .PCOut(PC), .MAROut(MAR), .MDROut(MDR), .IROut(IR));
regCC CCreg(.*, .CCIn(newCC), .BENIn(newBEN), .CCOut(CC), .BENOut(BEN));
reg_file GPR(.*, .SR1(SR1MUXOUT), .SR2(IR[2:0]), .DR(DRMUXOUT), .Din(databus));
ALU LC3ALU(.*, .A(SR1OUT), .B(SR2MUXOUT), .Out(ALUOut));

// Our SRAM and I/O controller (note, this plugs into MDR/MAR)

Mem2IO memory_subsystem(
    .*, .Reset(Reset), .ADDR(ADDR), .Switches(SW),
    .HEX0(hex_4[0][3:0]), .HEX1(hex_4[1][3:0]), .HEX2(hex_4[2][3:0]), .HEX3(hex_4[3][3:0]),
    .Data_from_CPU(MDR), .Data_to_CPU(MDR_In),
    .Data_from_SRAM(Data_from_SRAM), .Data_to_SRAM(Data_to_SRAM)
);

// State machine, you need to fill in the code here as well
ISDU state_controller(
	.*, .Reset(Reset), .Run(Run), .Continue(Continue),
	.Opcode(IR[15:12]), .IR_5(IR[5]), .IR_11(IR[11]),
   .Mem_OE(OE), .Mem_WE(WE)
);

// SRAM WE register
//logic SRAM_WE_In, SRAM_WE;
//// SRAM WE synchronizer
//always_ff @(posedge Clk or posedge Reset_ah)
//begin
//	if (Reset_ah) SRAM_WE <= 1'b1; //resets to 1
//	else 
//		SRAM_WE <= SRAM_WE_In;
//end

	
endmodule
